`include "uvm_macros.svh"
import uvm_pkg::*;

class seq_fifo_05 extends uvm_sequence #(apb_fifo_txn);
    `uvm_object_utils(seq_fifo_05)
    
    apb_fifo_vsqr vsqr;
    apb_fifo_seq wr_seq;
    apb_fifo_seq rd_seq;
    virtual apb_if vif;
    uvm_status_e status;
    uvm_reg_data_t read_val;
    
    function new(string name = "seq_fifo_05");
        super.new(name);
    endfunction

    /*
        TestID: FIFO_05
        Description: Write when full
    */
    task body();
        if (!$cast(vsqr, m_sequencer)) begin
            `uvm_fatal("FIFO_05", "Cannot cast m_sequencer to apb_fifo_vsqr")
        end

        // configure depth to 8
        vsqr.rgm.reg0.write(
            .status(status),
            .value(6'b00_0001),
            .parent(this),
            .path(UVM_FRONTDOOR)
        );

        for(int i=0;i<16;i++) begin
            wr_seq = apb_fifo_seq::type_id::create($sformatf("wr_0%d",i));
            wr_seq.op_type = FIFO_WRITE;
            wr_seq.gap_cycles = 0;
            wr_seq.start(vsqr.apb_sqr);
        end
    endtask
endclass