package apb_fifo_types_pkg;

  typedef enum {REG_CFG, REG_READ, FIFO_WRITE, FIFO_READ} apb_op_code;

endpackage
